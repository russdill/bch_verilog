`timescale 1ns / 1ps

`include "bch_defs.vh"

module sim #(
	parameter [`BCH_PARAM_SZ-1:0] P = `BCH_SANE,
	parameter OPTION = "SERIAL",
	parameter BITS = 1
) (
	input clk,
	input reset,
	input [`BCH_DATA_BITS(P)-1:0] data_in,
	input [`BCH_CODE_BITS(P)-1:0] error,
	input encode_start,
	output busy,
	output reg wrong = 0
);

`include "bch.vh"

localparam TCQ = 1;
localparam N = `BCH_N(P);
localparam E = `BCH_ECC_BITS(P);
localparam M = `BCH_M(P);
localparam T = `BCH_T(P);
localparam K = `BCH_K(P);
localparam B = `BCH_DATA_BITS(P);

reg [B-1:0] encode_buf = 0;
reg [E+B-1:0] flip_buf = 0;
reg [B-1:0] err_buf = 0;
reg last_data_valid = 0;

wire [BITS-1:0] encoded_data;
wire encoded_first;
wire encoded_last;
wire [BITS-1:0] decoder_in;
wire decode_busy;
wire encode_busy;
wire [`BCH_SYNDROMES_SZ(P)-1:0] syndromes;
wire syn_done;
wire err_start;
wire err_valid;
wire err;
wire key_busy;
wire errors_present;
wire [`BCH_ERR_SZ(P)-1:0] err_count;

assign busy = encode_busy;

localparam STACK_SZ = 6;

reg [STACK_SZ*`BCH_ERR_SZ(P)-1:0] err_count_stack = 0;
reg [STACK_SZ-1:0] err_present_stack = 0;
reg [STACK_SZ*`BCH_DATA_BITS(P)-1:0] err_stack = 0;

reg [log2(STACK_SZ)-1:0] wr_pos = 0;
reg [log2(STACK_SZ)-1:0] err_count_rd_pos = 0;
reg [log2(STACK_SZ)-1:0] err_present_rd_pos = 0;
reg [log2(STACK_SZ)-1:0] err_rd_pos = 0;

wire err_count_overflow = ((wr_pos + 1) % STACK_SZ) === err_count_rd_pos;
wire err_present_overflow = ((wr_pos + 1) % STACK_SZ) === err_present_rd_pos;
wire err_overflow = ((wr_pos + 1) % STACK_SZ) === err_rd_pos;

function integer bit_count;
	input [N-1:0] bits;
	integer count;
begin
	count = 0;
	while (bits) begin
		count = count + (bits[0] ? 1'b1 : 1'b0);
		bits = bits >> 1;
	end
	bit_count = count;
end
endfunction

always @(posedge clk) begin
	if (encode_start && !encode_busy && !decode_busy) begin
		err_stack[`BCH_DATA_BITS(P)*wr_pos+:`BCH_DATA_BITS(P)] <= #TCQ error;
		err_count_stack[`BCH_ERR_SZ(P)*wr_pos+:`BCH_ERR_SZ(P)] <= #TCQ bit_count(error);
		err_present_stack[wr_pos] <= #TCQ |error;
		wr_pos <= #TCQ (wr_pos + 1) % STACK_SZ;
	end

	if (!decode_busy) begin
		encode_buf <= #TCQ encode_start ? data_in : {{BITS{1'b0}}, encode_buf[`BCH_DATA_BITS(P)-1:BITS]};
		flip_buf   <= #TCQ encode_start ? error   : {{BITS{1'b0}}, flip_buf[`BCH_CODE_BITS(P)-1:BITS]};
	end
end

/* Generate code */
bch_encode #(P, BITS) u_bch_encode(
	.clk(clk),
	.start(encode_start),
	.data_in(encode_start ? data_in[BITS-1:0] : encode_buf[BITS*2-1:BITS]),
	.data_out(encoded_data),
	.first(encoded_first),
	.last(encoded_last),
	.accepted(!decode_busy),
	.busy(encode_busy)
);

assign decoder_in = encoded_data ^ flip_buf[BITS-1:0];

/* Process syndromes */
bch_syndrome #(P, BITS) u_bch_syndrome(
	.clk(clk),
	.start(encoded_first && !decode_busy),
	.busy(decode_busy),
	.data_in(decoder_in),
	.syndromes(syndromes),
	.done(syn_done),
	.accepted(syn_done && !key_busy)
);

/* Test for errors */
bch_errors_present #(P) u_errors(
	.start(syn_done && !key_busy),
	.syndromes(syndromes),
	.errors_present(errors_present)
);


wire err_present_wrong = syn_done && !key_busy && (errors_present !== err_present_stack[err_present_rd_pos]);

always @(posedge clk) begin
	if (syn_done && !key_busy)
		err_present_rd_pos = (err_present_rd_pos + 1) % STACK_SZ;
end

wire err_count_wrong;
if (OPTION == "SERIAL" || OPTION == "PARALLEL") begin : TMEC

	wire ch_start;
	wire ch_busy;
	wire [`BCH_SIGMA_SZ(P)-1:0] sigma;

	/* Solve key equation */
	if (OPTION == "SERIAL") begin : BMA_SERIAL
		bch_sigma_bma_serial #(P) u_bma (
			.clk(clk),
			.start(syn_done),
			.syndromes(syndromes),
			.sigma(sigma),
			.done(ch_start),
			.busy(key_busy),
			.accepted(!ch_busy),
			.err_count(err_count)
		);
	end else if (OPTION == "PARALLEL") begin : BMA_PARALLEL
		bch_sigma_bma_parallel #(P) u_bma (
			.clk(clk),
			.start(syn_done),
			.syndromes(syndromes),
			.sigma(sigma),
			.done(ch_start),
			.busy(key_busy),
			.accepted(!ch_busy),
			.err_count(err_count)
		);
	end

	assign err_count_wrong = ch_start && (err_count !== err_count_stack[err_count_rd_pos*`BCH_ERR_SZ(P)+:`BCH_ERR_SZ(P)]);
	always @(posedge clk) begin
		if (ch_start && !ch_busy)
			err_count_rd_pos <= #TCQ (err_count_rd_pos + 1) % STACK_SZ;
	end

	/* Locate errors */
	bch_error_tmec #(P) u_error_tmec(
		.clk(clk),
		.start(ch_start && !ch_busy),
		.busy(ch_busy),
		.accepted(1'b1),
		.sigma(sigma),
		.ready(err_start),
		.valid(err_valid),
		.err(err)
	);

end else begin : DEC

	/* Locate errors */
	bch_error_dec #(P) u_error_dec(
		.clk(clk),
		.start(syn_done),
		.busy(key_busy),
		.accepted(1'b1),
		.syndromes(syndromes),
		.ready(err_start),
		.valid(err_valid),
		.err(err),
		.err_count(err_count)
	);

	assign err_count_wrong = err_done && (err_count !== err_count_stack[err_count_rd_pos*`BCH_ERR_SZ(P)+:`BCH_ERR_SZ(P)]);
	always @(posedge clk) begin
		if (err_done)
			err_count_rd_pos <= #TCQ (err_count_rd_pos + 1) % STACK_SZ;
	end

end

wire err_done = last_err_valid && !err_valid;
reg last_err_valid = 0;

wire err_wrong = err_done && (err_buf !== err_stack[err_rd_pos*B+:B]);
wire new_wrong = err_count_overflow || err_overflow || err_present_wrong || err_count_wrong || err_wrong;

always @(posedge clk) begin
	last_err_valid <= #TCQ err_valid;
	if (err_start)
		err_buf <= #TCQ {err, {`BCH_DATA_BITS(P)-1{1'b0}}};
	else if (err_valid)
		err_buf <= #TCQ {err, err_buf[`BCH_DATA_BITS(P)-1:1]};

	if (err_done)
		err_rd_pos <= #TCQ (err_rd_pos + 1) % STACK_SZ;

	if (reset)
		wrong <= #TCQ 1'b0;
	else if (new_wrong)
		wrong <= #TCQ 1'b1;
end

endmodule
